`timescale 1ns / 1ps

module mystery_func(
    input a,
    input b,
    input c,
    input d,
    input e,
    input f,
    output y
    );
    
// Add internal wire definitons here.
//    wire int_sig1, int_sig2, int_sig3, int_sig4, int_sig5, int_sig6, int_sig7, int_sig8;
    
// Add Design Code here.
        
endmodule