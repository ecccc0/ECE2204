`timescale 1ns / 1ps

module three_inp_func(
    input a,
    input b,
    input c,
    output y
    );

// Add internal wire definitions here.
//    wire int_sig1, int_sig2, int_sig3, int_sig4;

// Add design code here.    
    
endmodule
